`define BRAM_CONFIG_SELECT  (2'h0)
`define BRAM_MOD_SELECT     (2'h1)
`define BRAM_TR_SELECT      (2'h2)
`define BRAM_SEQ_SELECT     (2'h3)

`define MOD_BRAM_ADDR_OFFSET_ADDR (14'h0006)
`define SEQ_BRAM_ADDR_OFFSET_ADDR (14'h0007)

`define SEQ_MODE_FOCI           (0)
`define SEQ_MODE_RAW_DUTY_PHASE (1)
