/*
 * File: mult.sv
 * Project: common
 * Created Date: 07/01/2022
 * Author: Shun Suzuki
 * -----
 * Last Modified: 07/01/2022
 * Modified By: Shun Suzuki (suzuki@hapis.k.u-tokyo.ac.jp)
 * -----
 * Copyright (c) 2022 Hapis Lab. All rights reserved.
 * 
 */

`timescale 1ns / 1ps
module mult#(
           parameter int WIDTH_A,
           parameter int WIDTH_B
       )(
           input var CLK,
           input var [WIDTH_A-1:0] A,
           input var [WIDTH_B-1:0] B,
           output var [WIDTH_A+WIDTH_B-1:0] P
       );

MULT_MACRO #(
               .DEVICE("7SERIES"),
               .LATENCY(3),
               .WIDTH_A(WIDTH_A),
               .WIDTH_B(WIDTH_B)
           ) MULT_MACRO_inst (
               .P(P),
               .A(A),
               .B(B),
               .CE(1'b1),
               .CLK(CLK),
               .RST()
           );

endmodule
